`timescale 1ns / 1ps
module I_cache(
    input wire
);