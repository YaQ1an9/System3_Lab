`ifndef I_STAGE_H
`define I_STAGE_H

parameter   IDLE = 2'b00,
            CompareTag = 2'b01,
            Allocate = 2'b

`endif