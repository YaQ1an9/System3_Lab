`ifndef I_STAGE_H
`define I_STAGE_H

parameter   IDLE = 3'b000,
            CompareTag = 3'b001,
            Allocate = 3'b10,
            WriteBack = 2'b11;

`endif