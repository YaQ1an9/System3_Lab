`ifndef I_STAGE_H
`define I_STAGE_H

parameter   

`endif