`ifndef STAGE_H
#