`timescale 1ns / 1ps

module MUX8T1_32(
    input [31:0] I0,
    input [31:0] I1,
    input [31:0] I2,
    input [31:0] I3,
    input [31:0] I4,
    input [31:0] I5,
    input [31:0] I6,
    input [31:0] I7,
    input [31:0] I8,
    input [1:0]Forward,
    input [1:0]src,
    output [31:0]o
    );
    always @(*)
    begin
    end
endmodule
