`timescale 1ns / 1ps
module I_cache(
    input wire clk,
    input wire rst,

    input [31:0] 
);