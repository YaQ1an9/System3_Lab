`ifndef STAGE_H
`