//`ifndef ALUOP_H
//`define ALUOP_H
parameter   ADD  = 4'b0000,
            SUB  = 4'b1000,
			SLL  = 4'b0001,
			SLT  = 4'b0010,
			SLTU = 4'b0011,
			XOR  = 4'b0100,
			SRL  = 4'b0101,
			SRA  = 4'b1101,
			OR   = 4'b0110,
			AND  = 4'b0111,
			NOP  = 4'b1111,
			CMP  = 4'b1010,
			CMP_U  = 4'b1001;
//`endif