`ifndef I_STAGE_H
`define I_STAGE_H

parameter   IDLE = 3'b000,
            CompareTag = 2'b01,
            Allocate = 2'b10,
            WriteBack = 2'b11;

`endif