`ifndef MEM_ACCESS_SIZE
`define MEM_ACCESS_SIZE
parameter Signed_Byte = 3'b000;
parameter Half_Word = 3'b001;
parameter Word = 3'b010;
parameter Unsigned_Byte = 3'b100;
parameter Double_Word = 3'b101;


`endif