`ifndef STAGE_H
`define STAGE_