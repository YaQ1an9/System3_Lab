//ifndef STAGE_H
#