`ifndef I_STAGE_H
`define I_STAGE_H

parameter   IDLE = 2'b00,
            

`endif