#ifndef STAGE_H
#