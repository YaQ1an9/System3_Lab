ifndef STAGE_H
#