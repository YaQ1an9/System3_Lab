`ifndef STAGE_H
`define STAGE_H

parameter   S_IDLE = 3'b0000,
            S_BACK = 3

`endif