`ifndef CSR_NUM
`define CSR_NUM
parameter sstatus = 12'h100;
parameter stvec = 12'h105;
parameter scause = 12'h142;
parameter satp = 12'h180;
parameter sepc = 12'h141;
parameter mstatus = 12'h300;
parameter mscratch = 12'h340;
parameter mepc = 12'h341;
parameter mcause = 12'h342;
parameter mtvec = 12'h305;
`endif