`ifndef STAGE_H
`define STAGE_H

parameter   

`e